-- THIS FILE IS OBSOLETE