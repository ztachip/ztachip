-- THIS FILE IS OBSOLETE. REPLACED WITH DDR_RX.VHD AND DDR_TX.VHD