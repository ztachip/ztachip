------------------------------------------------------------------------------
-- Copyright [2014] [Ztachip Technologies Inc]
--
-- Author: Vuong Nguyen
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
-- http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
------------------------------------------------------------------------------
----------
-- This module implements simple dual-port ram for Xilinx
----------

library std;
use std.standard.all;
LIBRARY ieee;
USE ieee.std_logic_1164.all;
use IEEE.numeric_std.all;
use work.ztachip_pkg.all;
Library xpm;
use xpm.vcomponents.all;

ENTITY DPRAM_DUAL_CLOCK IS
   GENERIC (
        numwords_a                      : NATURAL;
        numwords_b                      : NATURAL;
        widthad_a                       : NATURAL;
        widthad_b                       : NATURAL;
        width_a                         : NATURAL;
        width_b                         : NATURAL
    );
    PORT (
        address_a : IN STD_LOGIC_VECTOR (widthad_a-1 DOWNTO 0);
        clock_a   : IN STD_LOGIC;
        clock_b   : IN STD_LOGIC;
        data_a    : IN STD_LOGIC_VECTOR (width_a-1 DOWNTO 0);
        q_b       : OUT STD_LOGIC_VECTOR (width_b-1 DOWNTO 0);
        wren_a    : IN STD_LOGIC ;
        address_b : IN STD_LOGIC_VECTOR (widthad_b-1 DOWNTO 0)
    );
END DPRAM_DUAL_CLOCK;

architecture dpram_behaviour of DPRAM_DUAL_CLOCK is

SIGNAL byteena_a:std_logic_vector(0 downto 0);

begin

byteena_a(0) <= wren_a;

xpm_memory_sdpram_inst : xpm_memory_dpdistram
generic map (
    ADDR_WIDTH_A => widthad_a, -- DECIMAL
    ADDR_WIDTH_B => widthad_b, -- DECIMAL
    BYTE_WRITE_WIDTH_A => width_a, -- DECIMAL
    CLOCKING_MODE => "independent_clock", -- String
    MEMORY_INIT_FILE => "none", -- String
    MEMORY_INIT_PARAM => "0", -- String
    MEMORY_OPTIMIZATION => "true", -- String
    MEMORY_SIZE => numwords_a*width_a, -- DECIMAL
    MESSAGE_CONTROL => 0, -- DECIMAL
    READ_DATA_WIDTH_A => width_b, -- DECIMAL
    READ_DATA_WIDTH_B => width_b, -- DECIMAL
    READ_LATENCY_B => 1, -- DECIMAL
    READ_RESET_VALUE_B => "0", -- String
    RST_MODE_A => "SYNC", -- String
    RST_MODE_B => "SYNC", -- String
    SIM_ASSERT_CHK => 0, -- DECIMAL; 0=disable simulation messages, 1=enable simulation messages
    USE_EMBEDDED_CONSTRAINT => 1, -- DECIMAL
    USE_MEM_INIT => 1, -- DECIMAL
    USE_MEM_INIT_MMI => 0, -- DECIMAL
    WRITE_DATA_WIDTH_A => width_a
)
port map (
    doutb => q_b,         -- READ_DATA_WIDTH_B-bit output: Data output for port B read operations.
    addra => address_a,   -- ADDR_WIDTH_A-bit input: Address for port A write operations.
    addrb => address_b,   -- ADDR_WIDTH_B-bit input: Address for port B read operations.
    clka => clock_a,      -- 1-bit input: Clock signal for port A. Also clocks port B when
    clkb => clock_b,      -- 1-bit input: Clock signal for port B when parameter CLOCKING_MODE is
                          -- "independent_clock". Unused when parameter CLOCKING_MODE is
                          -- "common_clock".
    dina => data_a,       -- WRITE_DATA_WIDTH_A-bit input: Data input for port A write operations.
    ena => wren_a,        -- 1-bit input: Memory enable signal for port A. Must be high on clock
    enb => '1',           -- 1-bit input: Memory enable signal for port B. Must be high on clock
    regceb => '1',         -- 1-bit input: Clock Enable for the last register stage on the output
                           -- data path.
    rsta => '0',           -- 1-bit input: Reset signal for the final port B output register

    rstb => '0',           -- 1-bit input: Reset signal for the final port B output register
                           -- stage. Synchronously resets output port doutb to the value specified
                           -- by parameter READ_RESET_VALUE_B.
    wea => byteena_a,      -- WRITE_DATA_WIDTH_A/BYTE_WRITE_WIDTH_A-bit input: Write enable vector
                           -- for port A input data port dina. 1 bit wide when word-wide writes
                           -- are used. In byte-wide write configurations, each bit controls the
                           -- writing one byte of dina to address addra. For example, to
                           -- synchronously write only bits [15-8] of dina when WRITE_DATA_WIDTH_A
                           -- is 32, wea would be 4'b0010.
    regcea => '1'
);

end dpram_behaviour;
