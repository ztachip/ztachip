-- THIS FILE IS OBSOLETE ---